<!-- List of labels:
PREP Prepositions
PRNTONIC  *** not applicable ***
PRNSUBJ Subject form of personal pronouns
PRNOBJ Object form of personal pronouns
PRNPOS Possessive prounouns and determiners, incl. genitiv
PRNREF Reflexive/reciprocal pronouns
PRN any pronoun
ONLYPRN *** not applicable ***
CNJCOO Co-ordinating conjunction
CNJSUB Sub-ordinating conjunction
*** label for <sdef n="cnjadv" 	c="Adverbial conjunction"/> is missing ***

-->