<!-- List of labels:
PREP Prepositions

PRNTONIC  *** not applicable ***

PRNSUBJ Subject form of personal pronouns
PRNOBJ Object form of personal pronouns
PRNPOS Possessive prounouns and determiners, incl. genitiv
PRNREF Reflexive/reciprocal pronouns
PRN any pronoun

ONLYPRN *** not applicable ***

CNJCOO Co-ordinating conjunction
CNJSUB Sub-ordinating conjunction
CNJADV Adverbial conjunction

*** label for <sdef n="cnjadv" 	c="Adverbial conjunction"/> is missing ***

DETDEM Demonstrative pronoun
DETIND Indefinite determiner
DETDEF Definite determiner

DETPOS *** not in use: PRONPOS instead ***

DETORD Ordinal determiner (ordinal number)
DETQNT Quantifier
IJ Interjections

REL *** not applicable ***

NOMSDEF Definite noun
NOMSSING Noun in singular
NOMSPROPIS Proper noun
NOMSNEUTREUTRE Common gender or neuter *** not applicable ***
NOMSNEUTRE Noun, Neuter
NOMSUTRE Noun, Common gender (Utrum)

ADV Adverb

PREADV *** not applicable ***
ADVS *** not applicable ***
ADVPOS *** not applicable ***
CONJADV *** not applicable ***

ADJPLUR adjective in plural NEW
ADJ Adjective
NUM Numeral

NUMS *** not applicable ***
VBMODDA *** not applicable ***
VBMODPRET *** not applicable ***

VBMODINF Modal verb: infinitive
VBMODINFS Modal verb: infinitive + eg. active voice/passive voice
VBMODPRES Modal verb: presens
VBMODPRESS Modal verb: presens + eg. active voice/passive voice
VBMODPAST Modal verb: Past
VBMODPASTS Modal verb: Past + eg. active voice/passive voice
VBMODSUPN Modal verb: Supinum
VBMODPPRES Modal verb: Present participle
VBMODIMP Modal verb: Imperfekt NEW

VBAUXPRS *** not applicable ***
VBAUXDA *** not applicable ***
VBAUXPRET *** not applicable ***
VBAUXINF *** not applicable *** see VAUXINF etc!

VBSPRS *** not applicable ***
VBSDA *** not applicable ***
VBSPRET *** not applicable ***
VBSINF *** not applicable ***

VBLEXPRS Lexical (normal) verb: Present (presens)
VBLEXDA Lexical (normal) verb: Past
VBLEXPART Lexical (normal) verb: Past participle
VBLEXPPRES Lexical (normal) verb: Present participle
VBLEXINF Lexical (normal) verb: Infinitive
VBLEXSUPN Lexical (normal) verb: Supine (Supinum)
VBLEXSUPNS Lexical (normal) verb: Supine + eg. active voice
VBLEXPRET *** not defined ***

VBSERINF vbser (to be): infinitive
VBSERPAST vbser (to be): past
VBSERPRES vbser (to be): present
VBSERSUPN vbser (to be): Supine
VBSERPPRES vbser (to be): Present participle
VBSERPPRESS *** not applicable ***
VBSERIMP vbser (to be): imperfect NEW

VBHAVERPRES vbhaver (to have): present
VBHAVERPAST vbhaver (to have): past
VBHAVERPPRES vbhaver (to have): Present participle
VBHAVERINF vbhaver (to have): Infinitive
VBHAVERSUPN vbhaver (to have): Supine
VBHAVERPP vbhaver (to have): Past participl

VAUXINF auxilary verb: Infinitive
VAUXPRES auxilary verb: Present
VAUXPAST auxilary verb: Past
VAUXPASTS auxilary verb: *** Not used ***
VAUXSUPN auxilary verb: Supine
VAUXSUPNS auxilary verb: *** Not used ***

ADVH�R lemma 'h�r':  *** Not used ***

VBCLOSED all other vbser and vbhaver

VB all other lexical verbs (open)

-->









-->